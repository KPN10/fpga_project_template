module top (
    input logic i_clock
);

endmodule
